library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity four_bit_alu is
    Port (
	A : in STD_LOGIC_VECTOR (3 downto 0); 
	B : in STD_LOGIC_VECTOR (3 downto 0);
	Opcode : in STD_LOGIC_VECTOR (1 downto 0);
	Result : out STD_LOGIC_VECTOR (3 downto 0);
	Equal : out STD_LOGIC;
	Cout : out STD_LOGIC
    );
end four_bit_alu;

architecture Four_bit_alu is
signal temp_s: signed(4 downto 0) := (other => '0'); -- to hold temporary results, like your b register
begin
    process(A, B, Opcode)
    	begin
		case (Opcode) is
			when "00" =>
			temp_s <= signed('0' & A) + signed('0' & B);
			if (temp_s(4) /= temp(3)) then
				overflow <= '1';
			else
				overflow <= '0';
			end if;

			when "01" =>
			temp_s <= signed('0' & A) - signed('0' & B);
			if (temp_s(4) /= temp(3)) then
				overflow <= '1';
			else
				overflow <= '0';
			end if;

			when "10" =>
			temp_s <= A and B;

			when "11" =>
			temp_s <= A or B;
		end case;
	end process;
	process (A, B)
	begin
	     if (A = B) then
		Equal <= '1';
			else
				Equal <= '0';
	     end if;
	end process;
		Output <= STD_LOGIC_VECTOR(temp_s(3 downto 0));
		Overflow <= STD_LOGIC_VECTOR(temp_s(3));
    end process
end Four_bit_alu;

